module div(
	input [10000000:0]A,
	input [10000000:0]B,
	output [10000000:0]C
);

assign C = A/B;
endmodule
